
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h7c388cfe;
    ram_cell[       1] = 32'h0;  // 32'hd40c187d;
    ram_cell[       2] = 32'h0;  // 32'h6d9159c2;
    ram_cell[       3] = 32'h0;  // 32'ha0d7e4fa;
    ram_cell[       4] = 32'h0;  // 32'h1be35354;
    ram_cell[       5] = 32'h0;  // 32'h9b61c042;
    ram_cell[       6] = 32'h0;  // 32'h1fd79c26;
    ram_cell[       7] = 32'h0;  // 32'haaa00488;
    ram_cell[       8] = 32'h0;  // 32'h41c34993;
    ram_cell[       9] = 32'h0;  // 32'h7efcb998;
    ram_cell[      10] = 32'h0;  // 32'h9dd1b948;
    ram_cell[      11] = 32'h0;  // 32'h13c1cf11;
    ram_cell[      12] = 32'h0;  // 32'h78a849a5;
    ram_cell[      13] = 32'h0;  // 32'h622261e9;
    ram_cell[      14] = 32'h0;  // 32'h92f8c675;
    ram_cell[      15] = 32'h0;  // 32'heff37a14;
    ram_cell[      16] = 32'h0;  // 32'h48084789;
    ram_cell[      17] = 32'h0;  // 32'h3cab41f4;
    ram_cell[      18] = 32'h0;  // 32'hb0fcb42b;
    ram_cell[      19] = 32'h0;  // 32'h532b6f4e;
    ram_cell[      20] = 32'h0;  // 32'h4677d008;
    ram_cell[      21] = 32'h0;  // 32'hbb27c967;
    ram_cell[      22] = 32'h0;  // 32'h0a7597ec;
    ram_cell[      23] = 32'h0;  // 32'h88d9217d;
    ram_cell[      24] = 32'h0;  // 32'hd93343ef;
    ram_cell[      25] = 32'h0;  // 32'h6ef3eaa8;
    ram_cell[      26] = 32'h0;  // 32'hd35b3094;
    ram_cell[      27] = 32'h0;  // 32'h26684ffd;
    ram_cell[      28] = 32'h0;  // 32'hcb01a6de;
    ram_cell[      29] = 32'h0;  // 32'hf0dd7aef;
    ram_cell[      30] = 32'h0;  // 32'h89fdaff5;
    ram_cell[      31] = 32'h0;  // 32'h3c0aea56;
    ram_cell[      32] = 32'h0;  // 32'h6dfd5121;
    ram_cell[      33] = 32'h0;  // 32'hdea9eafe;
    ram_cell[      34] = 32'h0;  // 32'h2bd3671c;
    ram_cell[      35] = 32'h0;  // 32'hb1c62197;
    ram_cell[      36] = 32'h0;  // 32'hd7952074;
    ram_cell[      37] = 32'h0;  // 32'hef18ef55;
    ram_cell[      38] = 32'h0;  // 32'hc741d09e;
    ram_cell[      39] = 32'h0;  // 32'h2cf80705;
    ram_cell[      40] = 32'h0;  // 32'hd8fb3939;
    ram_cell[      41] = 32'h0;  // 32'h9d9528c7;
    ram_cell[      42] = 32'h0;  // 32'h72ce5022;
    ram_cell[      43] = 32'h0;  // 32'h53ef857a;
    ram_cell[      44] = 32'h0;  // 32'h6927bb4d;
    ram_cell[      45] = 32'h0;  // 32'h72965f99;
    ram_cell[      46] = 32'h0;  // 32'h32b921ea;
    ram_cell[      47] = 32'h0;  // 32'h24ed050e;
    ram_cell[      48] = 32'h0;  // 32'h38e7027a;
    ram_cell[      49] = 32'h0;  // 32'h76f7f678;
    ram_cell[      50] = 32'h0;  // 32'hfc95d4ee;
    ram_cell[      51] = 32'h0;  // 32'h469796a1;
    ram_cell[      52] = 32'h0;  // 32'h51404e34;
    ram_cell[      53] = 32'h0;  // 32'hf3501fcf;
    ram_cell[      54] = 32'h0;  // 32'hcb607297;
    ram_cell[      55] = 32'h0;  // 32'h9787e060;
    ram_cell[      56] = 32'h0;  // 32'hb5473ceb;
    ram_cell[      57] = 32'h0;  // 32'hecaeac9a;
    ram_cell[      58] = 32'h0;  // 32'h18d85c09;
    ram_cell[      59] = 32'h0;  // 32'h1e8f5986;
    ram_cell[      60] = 32'h0;  // 32'h57afef1a;
    ram_cell[      61] = 32'h0;  // 32'hc44adbc6;
    ram_cell[      62] = 32'h0;  // 32'hac1c3c06;
    ram_cell[      63] = 32'h0;  // 32'h6802587a;
    ram_cell[      64] = 32'h0;  // 32'h4a1b5213;
    ram_cell[      65] = 32'h0;  // 32'h771b7904;
    ram_cell[      66] = 32'h0;  // 32'h6481c28a;
    ram_cell[      67] = 32'h0;  // 32'hf8e06e89;
    ram_cell[      68] = 32'h0;  // 32'haf272b21;
    ram_cell[      69] = 32'h0;  // 32'h58dec468;
    ram_cell[      70] = 32'h0;  // 32'h6301fa62;
    ram_cell[      71] = 32'h0;  // 32'h283b5992;
    ram_cell[      72] = 32'h0;  // 32'hcd452e79;
    ram_cell[      73] = 32'h0;  // 32'h3f68edb9;
    ram_cell[      74] = 32'h0;  // 32'h25a95736;
    ram_cell[      75] = 32'h0;  // 32'hcd5351ac;
    ram_cell[      76] = 32'h0;  // 32'hf0dcd14a;
    ram_cell[      77] = 32'h0;  // 32'hd6075ecc;
    ram_cell[      78] = 32'h0;  // 32'h8eb336cf;
    ram_cell[      79] = 32'h0;  // 32'hdba4d8d8;
    ram_cell[      80] = 32'h0;  // 32'hd782bd5f;
    ram_cell[      81] = 32'h0;  // 32'haf6d0f8d;
    ram_cell[      82] = 32'h0;  // 32'hdc4d08d7;
    ram_cell[      83] = 32'h0;  // 32'h9bb943e3;
    ram_cell[      84] = 32'h0;  // 32'h3f1b6e42;
    ram_cell[      85] = 32'h0;  // 32'h02322a27;
    ram_cell[      86] = 32'h0;  // 32'h3a793aac;
    ram_cell[      87] = 32'h0;  // 32'hd3701bf4;
    ram_cell[      88] = 32'h0;  // 32'h98288fd6;
    ram_cell[      89] = 32'h0;  // 32'h9986fcd9;
    ram_cell[      90] = 32'h0;  // 32'h82af5ca9;
    ram_cell[      91] = 32'h0;  // 32'hbf0cfef0;
    ram_cell[      92] = 32'h0;  // 32'h801c510e;
    ram_cell[      93] = 32'h0;  // 32'ha3c3a707;
    ram_cell[      94] = 32'h0;  // 32'he020e3e7;
    ram_cell[      95] = 32'h0;  // 32'h719d4aa1;
    ram_cell[      96] = 32'h0;  // 32'h6d6d596f;
    ram_cell[      97] = 32'h0;  // 32'h44e42793;
    ram_cell[      98] = 32'h0;  // 32'hfa77538e;
    ram_cell[      99] = 32'h0;  // 32'h0f1fbe77;
    ram_cell[     100] = 32'h0;  // 32'hccde8c0e;
    ram_cell[     101] = 32'h0;  // 32'h9a864628;
    ram_cell[     102] = 32'h0;  // 32'h23847f2a;
    ram_cell[     103] = 32'h0;  // 32'hf76b851d;
    ram_cell[     104] = 32'h0;  // 32'h7670584f;
    ram_cell[     105] = 32'h0;  // 32'hcf2684d0;
    ram_cell[     106] = 32'h0;  // 32'h61ef2f02;
    ram_cell[     107] = 32'h0;  // 32'h8701b3c4;
    ram_cell[     108] = 32'h0;  // 32'hf2c0e0e7;
    ram_cell[     109] = 32'h0;  // 32'h2f8e33ba;
    ram_cell[     110] = 32'h0;  // 32'he77d5431;
    ram_cell[     111] = 32'h0;  // 32'hc34befee;
    ram_cell[     112] = 32'h0;  // 32'ha689b610;
    ram_cell[     113] = 32'h0;  // 32'h2b65bca8;
    ram_cell[     114] = 32'h0;  // 32'hb3041e56;
    ram_cell[     115] = 32'h0;  // 32'h3ec6b42a;
    ram_cell[     116] = 32'h0;  // 32'h033dd47f;
    ram_cell[     117] = 32'h0;  // 32'h3f6738ce;
    ram_cell[     118] = 32'h0;  // 32'hff954791;
    ram_cell[     119] = 32'h0;  // 32'ha92e8a1b;
    ram_cell[     120] = 32'h0;  // 32'h6efccba8;
    ram_cell[     121] = 32'h0;  // 32'hddcb57df;
    ram_cell[     122] = 32'h0;  // 32'h07837397;
    ram_cell[     123] = 32'h0;  // 32'hd19674f8;
    ram_cell[     124] = 32'h0;  // 32'h6d04c718;
    ram_cell[     125] = 32'h0;  // 32'h857341b1;
    ram_cell[     126] = 32'h0;  // 32'habd0a3da;
    ram_cell[     127] = 32'h0;  // 32'h035e70e9;
    ram_cell[     128] = 32'h0;  // 32'hae579a8e;
    ram_cell[     129] = 32'h0;  // 32'hbfd7028d;
    ram_cell[     130] = 32'h0;  // 32'h252813ff;
    ram_cell[     131] = 32'h0;  // 32'h925f28bc;
    ram_cell[     132] = 32'h0;  // 32'h483a60f0;
    ram_cell[     133] = 32'h0;  // 32'h12a60d88;
    ram_cell[     134] = 32'h0;  // 32'ha37bfabc;
    ram_cell[     135] = 32'h0;  // 32'hfda9a6e3;
    ram_cell[     136] = 32'h0;  // 32'h6df258d0;
    ram_cell[     137] = 32'h0;  // 32'h75b8a7b2;
    ram_cell[     138] = 32'h0;  // 32'h3a126919;
    ram_cell[     139] = 32'h0;  // 32'h856eb7b2;
    ram_cell[     140] = 32'h0;  // 32'hab14ff9e;
    ram_cell[     141] = 32'h0;  // 32'h39ee5693;
    ram_cell[     142] = 32'h0;  // 32'hc31c7963;
    ram_cell[     143] = 32'h0;  // 32'h27d26e3d;
    ram_cell[     144] = 32'h0;  // 32'h8610ff66;
    ram_cell[     145] = 32'h0;  // 32'ha2858afc;
    ram_cell[     146] = 32'h0;  // 32'h5c4f20c9;
    ram_cell[     147] = 32'h0;  // 32'hb0c2fa77;
    ram_cell[     148] = 32'h0;  // 32'h0450dc2f;
    ram_cell[     149] = 32'h0;  // 32'h1d115e83;
    ram_cell[     150] = 32'h0;  // 32'h5ebf4cb2;
    ram_cell[     151] = 32'h0;  // 32'hc2ad5d8c;
    ram_cell[     152] = 32'h0;  // 32'hac5d1902;
    ram_cell[     153] = 32'h0;  // 32'hf274a9e4;
    ram_cell[     154] = 32'h0;  // 32'h20ad9207;
    ram_cell[     155] = 32'h0;  // 32'h969e6c61;
    ram_cell[     156] = 32'h0;  // 32'h9e05f8bf;
    ram_cell[     157] = 32'h0;  // 32'h0138f5fd;
    ram_cell[     158] = 32'h0;  // 32'h24c6139f;
    ram_cell[     159] = 32'h0;  // 32'h7234403f;
    ram_cell[     160] = 32'h0;  // 32'h1ef9df8b;
    ram_cell[     161] = 32'h0;  // 32'h8fa956a0;
    ram_cell[     162] = 32'h0;  // 32'h0597df8c;
    ram_cell[     163] = 32'h0;  // 32'h79f20c9f;
    ram_cell[     164] = 32'h0;  // 32'h1d17e195;
    ram_cell[     165] = 32'h0;  // 32'h1b75592c;
    ram_cell[     166] = 32'h0;  // 32'h762cb177;
    ram_cell[     167] = 32'h0;  // 32'h8a57ff47;
    ram_cell[     168] = 32'h0;  // 32'hbd227839;
    ram_cell[     169] = 32'h0;  // 32'h6b39a5a2;
    ram_cell[     170] = 32'h0;  // 32'h1a60ee82;
    ram_cell[     171] = 32'h0;  // 32'h7bfcb1e5;
    ram_cell[     172] = 32'h0;  // 32'h3fe51269;
    ram_cell[     173] = 32'h0;  // 32'h7d796181;
    ram_cell[     174] = 32'h0;  // 32'hc5217d53;
    ram_cell[     175] = 32'h0;  // 32'hb1ac1ff2;
    ram_cell[     176] = 32'h0;  // 32'h99c8f295;
    ram_cell[     177] = 32'h0;  // 32'h346042f2;
    ram_cell[     178] = 32'h0;  // 32'hbf4c9529;
    ram_cell[     179] = 32'h0;  // 32'he299d93d;
    ram_cell[     180] = 32'h0;  // 32'h2483adfa;
    ram_cell[     181] = 32'h0;  // 32'h02c627c6;
    ram_cell[     182] = 32'h0;  // 32'hf00dd3c5;
    ram_cell[     183] = 32'h0;  // 32'he49dade3;
    ram_cell[     184] = 32'h0;  // 32'h539aaef9;
    ram_cell[     185] = 32'h0;  // 32'hbe461053;
    ram_cell[     186] = 32'h0;  // 32'h170d9bfb;
    ram_cell[     187] = 32'h0;  // 32'h2ab13708;
    ram_cell[     188] = 32'h0;  // 32'hc04953f5;
    ram_cell[     189] = 32'h0;  // 32'h7c1d0f0e;
    ram_cell[     190] = 32'h0;  // 32'hacec0e51;
    ram_cell[     191] = 32'h0;  // 32'h147173a3;
    ram_cell[     192] = 32'h0;  // 32'h138dfc47;
    ram_cell[     193] = 32'h0;  // 32'hdef74912;
    ram_cell[     194] = 32'h0;  // 32'he024086f;
    ram_cell[     195] = 32'h0;  // 32'h63b2098a;
    ram_cell[     196] = 32'h0;  // 32'h5109fbbb;
    ram_cell[     197] = 32'h0;  // 32'hcc4e68fc;
    ram_cell[     198] = 32'h0;  // 32'h6cc9c11a;
    ram_cell[     199] = 32'h0;  // 32'h59be7229;
    ram_cell[     200] = 32'h0;  // 32'h7de19b62;
    ram_cell[     201] = 32'h0;  // 32'hfb0bc2a3;
    ram_cell[     202] = 32'h0;  // 32'h5e0d6540;
    ram_cell[     203] = 32'h0;  // 32'h4b66159d;
    ram_cell[     204] = 32'h0;  // 32'h427489a8;
    ram_cell[     205] = 32'h0;  // 32'h23092b2b;
    ram_cell[     206] = 32'h0;  // 32'hc0ee6f42;
    ram_cell[     207] = 32'h0;  // 32'hea06eca8;
    ram_cell[     208] = 32'h0;  // 32'ha31b42aa;
    ram_cell[     209] = 32'h0;  // 32'hebb8f88b;
    ram_cell[     210] = 32'h0;  // 32'heea9eda4;
    ram_cell[     211] = 32'h0;  // 32'h97a71385;
    ram_cell[     212] = 32'h0;  // 32'hea4b2a73;
    ram_cell[     213] = 32'h0;  // 32'h2e2bfa5a;
    ram_cell[     214] = 32'h0;  // 32'h464363d4;
    ram_cell[     215] = 32'h0;  // 32'h55dcb901;
    ram_cell[     216] = 32'h0;  // 32'h71478333;
    ram_cell[     217] = 32'h0;  // 32'h4b71def8;
    ram_cell[     218] = 32'h0;  // 32'h1b394fd4;
    ram_cell[     219] = 32'h0;  // 32'h4a30eb45;
    ram_cell[     220] = 32'h0;  // 32'h2e56d2bf;
    ram_cell[     221] = 32'h0;  // 32'hac46e6f7;
    ram_cell[     222] = 32'h0;  // 32'h27730fb5;
    ram_cell[     223] = 32'h0;  // 32'hdeea63b4;
    ram_cell[     224] = 32'h0;  // 32'ha8fecae4;
    ram_cell[     225] = 32'h0;  // 32'h2d52f819;
    ram_cell[     226] = 32'h0;  // 32'h714275f3;
    ram_cell[     227] = 32'h0;  // 32'h76f87cd9;
    ram_cell[     228] = 32'h0;  // 32'h40167c4a;
    ram_cell[     229] = 32'h0;  // 32'he09c2706;
    ram_cell[     230] = 32'h0;  // 32'h63bbb300;
    ram_cell[     231] = 32'h0;  // 32'h1ff997fd;
    ram_cell[     232] = 32'h0;  // 32'h0c5d1389;
    ram_cell[     233] = 32'h0;  // 32'h6e6ae6e8;
    ram_cell[     234] = 32'h0;  // 32'he86720a2;
    ram_cell[     235] = 32'h0;  // 32'h722b776c;
    ram_cell[     236] = 32'h0;  // 32'hf7246511;
    ram_cell[     237] = 32'h0;  // 32'h9094e924;
    ram_cell[     238] = 32'h0;  // 32'h4584b87a;
    ram_cell[     239] = 32'h0;  // 32'h17ba3352;
    ram_cell[     240] = 32'h0;  // 32'h0f3a8c80;
    ram_cell[     241] = 32'h0;  // 32'h668e082e;
    ram_cell[     242] = 32'h0;  // 32'h5a533454;
    ram_cell[     243] = 32'h0;  // 32'he552bd3d;
    ram_cell[     244] = 32'h0;  // 32'h00d93d30;
    ram_cell[     245] = 32'h0;  // 32'h0fe30418;
    ram_cell[     246] = 32'h0;  // 32'h6933199e;
    ram_cell[     247] = 32'h0;  // 32'h5a69ea1c;
    ram_cell[     248] = 32'h0;  // 32'h0e3556c2;
    ram_cell[     249] = 32'h0;  // 32'hff1ff529;
    ram_cell[     250] = 32'h0;  // 32'h30857c05;
    ram_cell[     251] = 32'h0;  // 32'h4abbce36;
    ram_cell[     252] = 32'h0;  // 32'hfe4e88aa;
    ram_cell[     253] = 32'h0;  // 32'he7a81685;
    ram_cell[     254] = 32'h0;  // 32'h7ef94d31;
    ram_cell[     255] = 32'h0;  // 32'hd1f57f27;
    // src matrix A
    ram_cell[     256] = 32'h80b57d35;
    ram_cell[     257] = 32'he1961a66;
    ram_cell[     258] = 32'h77fbd5c5;
    ram_cell[     259] = 32'h0919e6c2;
    ram_cell[     260] = 32'h92f3e357;
    ram_cell[     261] = 32'h07ff733a;
    ram_cell[     262] = 32'hf3cc38d4;
    ram_cell[     263] = 32'h71ea22a1;
    ram_cell[     264] = 32'h15329e1a;
    ram_cell[     265] = 32'hcc5c1ac0;
    ram_cell[     266] = 32'h9ff7ce6e;
    ram_cell[     267] = 32'h2b61dda1;
    ram_cell[     268] = 32'h4c7fe3b7;
    ram_cell[     269] = 32'h0157f8c2;
    ram_cell[     270] = 32'h2538cc2e;
    ram_cell[     271] = 32'h0b31c798;
    ram_cell[     272] = 32'hfdcfe03d;
    ram_cell[     273] = 32'h5175ae20;
    ram_cell[     274] = 32'h0fd0e6e4;
    ram_cell[     275] = 32'hb94d8dd6;
    ram_cell[     276] = 32'hba1dda15;
    ram_cell[     277] = 32'h31f1d9de;
    ram_cell[     278] = 32'h14b738dc;
    ram_cell[     279] = 32'h80910c80;
    ram_cell[     280] = 32'h99953d0a;
    ram_cell[     281] = 32'h129db500;
    ram_cell[     282] = 32'hd1277482;
    ram_cell[     283] = 32'hdfc90939;
    ram_cell[     284] = 32'h682f036e;
    ram_cell[     285] = 32'hec031133;
    ram_cell[     286] = 32'hd398bde4;
    ram_cell[     287] = 32'h435aa323;
    ram_cell[     288] = 32'h54909f35;
    ram_cell[     289] = 32'hb0eb62ae;
    ram_cell[     290] = 32'h8a9bbc04;
    ram_cell[     291] = 32'h60f0552a;
    ram_cell[     292] = 32'hfae5835b;
    ram_cell[     293] = 32'h1446fa0d;
    ram_cell[     294] = 32'hc40607e2;
    ram_cell[     295] = 32'h669eea80;
    ram_cell[     296] = 32'h88520f2c;
    ram_cell[     297] = 32'h1208d74a;
    ram_cell[     298] = 32'ha09e2760;
    ram_cell[     299] = 32'ha23b772b;
    ram_cell[     300] = 32'h42f81673;
    ram_cell[     301] = 32'hde5ef94d;
    ram_cell[     302] = 32'h9a96cff8;
    ram_cell[     303] = 32'h455383bb;
    ram_cell[     304] = 32'h9e4616c7;
    ram_cell[     305] = 32'hb1df28ff;
    ram_cell[     306] = 32'h96df65e4;
    ram_cell[     307] = 32'h17c11afe;
    ram_cell[     308] = 32'hd70b3d67;
    ram_cell[     309] = 32'he5bba9c0;
    ram_cell[     310] = 32'h282c7ffb;
    ram_cell[     311] = 32'h84fab9b8;
    ram_cell[     312] = 32'h571d9ea8;
    ram_cell[     313] = 32'h6ff294d5;
    ram_cell[     314] = 32'h9e7c42d0;
    ram_cell[     315] = 32'ha9248c15;
    ram_cell[     316] = 32'h55acc846;
    ram_cell[     317] = 32'hba78929b;
    ram_cell[     318] = 32'h5303bf1a;
    ram_cell[     319] = 32'h21b862a8;
    ram_cell[     320] = 32'h88128109;
    ram_cell[     321] = 32'h62f412cd;
    ram_cell[     322] = 32'hc1a51716;
    ram_cell[     323] = 32'h456e25cf;
    ram_cell[     324] = 32'hb440c138;
    ram_cell[     325] = 32'hfd416031;
    ram_cell[     326] = 32'hbc24d199;
    ram_cell[     327] = 32'h6a2057b5;
    ram_cell[     328] = 32'h6879b084;
    ram_cell[     329] = 32'ha850c35e;
    ram_cell[     330] = 32'h93e1b959;
    ram_cell[     331] = 32'h32a02329;
    ram_cell[     332] = 32'h1eb6cacf;
    ram_cell[     333] = 32'h2e092e7b;
    ram_cell[     334] = 32'hf9bcd157;
    ram_cell[     335] = 32'ha4138bed;
    ram_cell[     336] = 32'h21d0c6e7;
    ram_cell[     337] = 32'hed0427cb;
    ram_cell[     338] = 32'h51c95098;
    ram_cell[     339] = 32'h59e2b9ce;
    ram_cell[     340] = 32'h0f516b35;
    ram_cell[     341] = 32'he37e7e67;
    ram_cell[     342] = 32'h02e0dc44;
    ram_cell[     343] = 32'h49ff2730;
    ram_cell[     344] = 32'h1ed28344;
    ram_cell[     345] = 32'hdb6f671c;
    ram_cell[     346] = 32'hffef362d;
    ram_cell[     347] = 32'h7959a49c;
    ram_cell[     348] = 32'h6ba8aeae;
    ram_cell[     349] = 32'hdfd6268b;
    ram_cell[     350] = 32'h0a727613;
    ram_cell[     351] = 32'h609a4a35;
    ram_cell[     352] = 32'h99fcc863;
    ram_cell[     353] = 32'hc32f9377;
    ram_cell[     354] = 32'h618a70c4;
    ram_cell[     355] = 32'h9c826f54;
    ram_cell[     356] = 32'hdb360540;
    ram_cell[     357] = 32'h501fe914;
    ram_cell[     358] = 32'h91e4d530;
    ram_cell[     359] = 32'h5a112a01;
    ram_cell[     360] = 32'h661e77c2;
    ram_cell[     361] = 32'h592269bd;
    ram_cell[     362] = 32'h278a5112;
    ram_cell[     363] = 32'hd89816cd;
    ram_cell[     364] = 32'h4ca99b80;
    ram_cell[     365] = 32'h965a14fc;
    ram_cell[     366] = 32'h4cd419e2;
    ram_cell[     367] = 32'h49ffd0d0;
    ram_cell[     368] = 32'h808886c4;
    ram_cell[     369] = 32'hed27d56b;
    ram_cell[     370] = 32'hda4973cd;
    ram_cell[     371] = 32'h96cdbdde;
    ram_cell[     372] = 32'h87d6e443;
    ram_cell[     373] = 32'h5ffed3e2;
    ram_cell[     374] = 32'h9002b9e4;
    ram_cell[     375] = 32'h0f38e46c;
    ram_cell[     376] = 32'h76c32faf;
    ram_cell[     377] = 32'hb4299e43;
    ram_cell[     378] = 32'h123b822b;
    ram_cell[     379] = 32'he6de8c0f;
    ram_cell[     380] = 32'h9ed68a68;
    ram_cell[     381] = 32'h70a368c7;
    ram_cell[     382] = 32'h7bfcb1a5;
    ram_cell[     383] = 32'h6e608c2c;
    ram_cell[     384] = 32'h5fa82128;
    ram_cell[     385] = 32'h5a8c146f;
    ram_cell[     386] = 32'hb0d8a063;
    ram_cell[     387] = 32'hc3ec3f02;
    ram_cell[     388] = 32'h900e8ef7;
    ram_cell[     389] = 32'ha918fad2;
    ram_cell[     390] = 32'h77990c7a;
    ram_cell[     391] = 32'hcaaed5d1;
    ram_cell[     392] = 32'h3e855480;
    ram_cell[     393] = 32'h6da2e2a3;
    ram_cell[     394] = 32'haa857b25;
    ram_cell[     395] = 32'h49a281ec;
    ram_cell[     396] = 32'h6a50be4b;
    ram_cell[     397] = 32'h282fd474;
    ram_cell[     398] = 32'hafa17c2f;
    ram_cell[     399] = 32'h07e72abf;
    ram_cell[     400] = 32'h55ee398e;
    ram_cell[     401] = 32'h3cdfff0d;
    ram_cell[     402] = 32'h9e48843a;
    ram_cell[     403] = 32'h180a89e6;
    ram_cell[     404] = 32'h953e813b;
    ram_cell[     405] = 32'hd33aa881;
    ram_cell[     406] = 32'hd7e8755f;
    ram_cell[     407] = 32'h0edb9467;
    ram_cell[     408] = 32'h34cfdb28;
    ram_cell[     409] = 32'h43beda38;
    ram_cell[     410] = 32'hb430bc6a;
    ram_cell[     411] = 32'he7319f2f;
    ram_cell[     412] = 32'hfe2ba5ed;
    ram_cell[     413] = 32'h7216e111;
    ram_cell[     414] = 32'h7db13322;
    ram_cell[     415] = 32'hc4bdecfa;
    ram_cell[     416] = 32'hcbfee1e5;
    ram_cell[     417] = 32'hc32a1ff3;
    ram_cell[     418] = 32'hc9720430;
    ram_cell[     419] = 32'hac6201f6;
    ram_cell[     420] = 32'h7121684f;
    ram_cell[     421] = 32'h015f802c;
    ram_cell[     422] = 32'h0c71405f;
    ram_cell[     423] = 32'h6d5d3173;
    ram_cell[     424] = 32'h2a6bfc7f;
    ram_cell[     425] = 32'hca51716f;
    ram_cell[     426] = 32'h1975984f;
    ram_cell[     427] = 32'h4c550b84;
    ram_cell[     428] = 32'hf8000173;
    ram_cell[     429] = 32'ha8909312;
    ram_cell[     430] = 32'hdced4e0e;
    ram_cell[     431] = 32'hd2d6d64f;
    ram_cell[     432] = 32'h1ca22bc8;
    ram_cell[     433] = 32'he37e5b1b;
    ram_cell[     434] = 32'he62b43e3;
    ram_cell[     435] = 32'hf253c63f;
    ram_cell[     436] = 32'hee72c422;
    ram_cell[     437] = 32'h6a39f5eb;
    ram_cell[     438] = 32'h1e5eb21e;
    ram_cell[     439] = 32'h1a805303;
    ram_cell[     440] = 32'h37521902;
    ram_cell[     441] = 32'h32a62e3d;
    ram_cell[     442] = 32'h84970fce;
    ram_cell[     443] = 32'h0bd16eed;
    ram_cell[     444] = 32'h86f23c5e;
    ram_cell[     445] = 32'h0b11d499;
    ram_cell[     446] = 32'hd282cb7c;
    ram_cell[     447] = 32'h150a288f;
    ram_cell[     448] = 32'h2095fe1a;
    ram_cell[     449] = 32'hb5c7d875;
    ram_cell[     450] = 32'ha1e7e1a2;
    ram_cell[     451] = 32'h8277183b;
    ram_cell[     452] = 32'h4b31bbfa;
    ram_cell[     453] = 32'had899f4f;
    ram_cell[     454] = 32'h3495f224;
    ram_cell[     455] = 32'h5883f63b;
    ram_cell[     456] = 32'hb54f44fa;
    ram_cell[     457] = 32'h131614f5;
    ram_cell[     458] = 32'h0b123ac0;
    ram_cell[     459] = 32'hd53c7c68;
    ram_cell[     460] = 32'ha91df7f8;
    ram_cell[     461] = 32'h58d33ecd;
    ram_cell[     462] = 32'h634cfcf1;
    ram_cell[     463] = 32'h590574a4;
    ram_cell[     464] = 32'h8378be41;
    ram_cell[     465] = 32'h63257a70;
    ram_cell[     466] = 32'h48e6ed4a;
    ram_cell[     467] = 32'hfe6b6aa5;
    ram_cell[     468] = 32'h0bc659a3;
    ram_cell[     469] = 32'h92bab533;
    ram_cell[     470] = 32'h0dbba0a4;
    ram_cell[     471] = 32'h6fc5cd9a;
    ram_cell[     472] = 32'hadfdd916;
    ram_cell[     473] = 32'h9f4d569e;
    ram_cell[     474] = 32'h21225e00;
    ram_cell[     475] = 32'h806069a8;
    ram_cell[     476] = 32'h6c0e922c;
    ram_cell[     477] = 32'hd1f95b71;
    ram_cell[     478] = 32'h564850c9;
    ram_cell[     479] = 32'h88c55a20;
    ram_cell[     480] = 32'hf72ab36a;
    ram_cell[     481] = 32'h8bf04a4f;
    ram_cell[     482] = 32'hdd5fe196;
    ram_cell[     483] = 32'h4803a773;
    ram_cell[     484] = 32'h853cac63;
    ram_cell[     485] = 32'h089cea29;
    ram_cell[     486] = 32'hb05d287a;
    ram_cell[     487] = 32'h17802686;
    ram_cell[     488] = 32'h79863079;
    ram_cell[     489] = 32'h82d64ac1;
    ram_cell[     490] = 32'haa84feb2;
    ram_cell[     491] = 32'h4d5ca76f;
    ram_cell[     492] = 32'h20dd890c;
    ram_cell[     493] = 32'hf699864a;
    ram_cell[     494] = 32'hb239fd67;
    ram_cell[     495] = 32'h12a23d85;
    ram_cell[     496] = 32'hc235b011;
    ram_cell[     497] = 32'h8a002096;
    ram_cell[     498] = 32'h26671711;
    ram_cell[     499] = 32'h0a327229;
    ram_cell[     500] = 32'h405ea51b;
    ram_cell[     501] = 32'h50c1a251;
    ram_cell[     502] = 32'hffe65ff3;
    ram_cell[     503] = 32'h5d672e4a;
    ram_cell[     504] = 32'h07f285da;
    ram_cell[     505] = 32'ha7d38deb;
    ram_cell[     506] = 32'hec3734dc;
    ram_cell[     507] = 32'hdab84df7;
    ram_cell[     508] = 32'h6504b5ab;
    ram_cell[     509] = 32'h0a3dfda9;
    ram_cell[     510] = 32'h27834ea3;
    ram_cell[     511] = 32'h56a82b19;
    // src matrix B
    ram_cell[     512] = 32'hb128f9d7;
    ram_cell[     513] = 32'h45bd536b;
    ram_cell[     514] = 32'hdfa7bbe9;
    ram_cell[     515] = 32'h6a8d4f6f;
    ram_cell[     516] = 32'h083e7abf;
    ram_cell[     517] = 32'ha03115b9;
    ram_cell[     518] = 32'hd0e55ddf;
    ram_cell[     519] = 32'hdf8639bb;
    ram_cell[     520] = 32'hb9b9b0f3;
    ram_cell[     521] = 32'h04ba323d;
    ram_cell[     522] = 32'hefdb3e69;
    ram_cell[     523] = 32'h97eaca07;
    ram_cell[     524] = 32'h37f057ba;
    ram_cell[     525] = 32'h3ac48c6a;
    ram_cell[     526] = 32'hda985cdc;
    ram_cell[     527] = 32'h21778928;
    ram_cell[     528] = 32'hc3175ac2;
    ram_cell[     529] = 32'h9d47f540;
    ram_cell[     530] = 32'h48505ca0;
    ram_cell[     531] = 32'h1d5a51e2;
    ram_cell[     532] = 32'hff1db241;
    ram_cell[     533] = 32'h07fae9b2;
    ram_cell[     534] = 32'h6620dfda;
    ram_cell[     535] = 32'he0084ab7;
    ram_cell[     536] = 32'h9ad1a4e7;
    ram_cell[     537] = 32'h59c7223f;
    ram_cell[     538] = 32'h9d0cdf2b;
    ram_cell[     539] = 32'hd2b9a1af;
    ram_cell[     540] = 32'h9ca91122;
    ram_cell[     541] = 32'h9ec97ff2;
    ram_cell[     542] = 32'h514b2627;
    ram_cell[     543] = 32'h827371a0;
    ram_cell[     544] = 32'ha8e9be1e;
    ram_cell[     545] = 32'h7d40a993;
    ram_cell[     546] = 32'h39cb8725;
    ram_cell[     547] = 32'hb767a59e;
    ram_cell[     548] = 32'hd4ffc718;
    ram_cell[     549] = 32'h4771bb42;
    ram_cell[     550] = 32'hc7ef62f6;
    ram_cell[     551] = 32'h6c17453a;
    ram_cell[     552] = 32'hfc6d1129;
    ram_cell[     553] = 32'h37f190bd;
    ram_cell[     554] = 32'hf335f911;
    ram_cell[     555] = 32'heece4dcc;
    ram_cell[     556] = 32'hefa7d84a;
    ram_cell[     557] = 32'h89e8cf46;
    ram_cell[     558] = 32'hd8d91db7;
    ram_cell[     559] = 32'h1a82032d;
    ram_cell[     560] = 32'hde0d7eab;
    ram_cell[     561] = 32'hc8cff24d;
    ram_cell[     562] = 32'h832e91df;
    ram_cell[     563] = 32'h28143450;
    ram_cell[     564] = 32'h6d651e16;
    ram_cell[     565] = 32'h4698e279;
    ram_cell[     566] = 32'hd84fdd3b;
    ram_cell[     567] = 32'hb238323f;
    ram_cell[     568] = 32'h496737b0;
    ram_cell[     569] = 32'he34265f3;
    ram_cell[     570] = 32'hc56c389b;
    ram_cell[     571] = 32'hc11197ca;
    ram_cell[     572] = 32'hc1a4eab9;
    ram_cell[     573] = 32'hcb139645;
    ram_cell[     574] = 32'hd904aec0;
    ram_cell[     575] = 32'h5a46e049;
    ram_cell[     576] = 32'hd8e258b1;
    ram_cell[     577] = 32'hfbfde30f;
    ram_cell[     578] = 32'hfd18128b;
    ram_cell[     579] = 32'h5ac15888;
    ram_cell[     580] = 32'h31c8a2ac;
    ram_cell[     581] = 32'h936c52da;
    ram_cell[     582] = 32'ha16f0883;
    ram_cell[     583] = 32'h0a0fc2e7;
    ram_cell[     584] = 32'hd88627b7;
    ram_cell[     585] = 32'hb4bfc8c7;
    ram_cell[     586] = 32'hffca401b;
    ram_cell[     587] = 32'hff3e3ab7;
    ram_cell[     588] = 32'h4cd1c9bd;
    ram_cell[     589] = 32'h7b721f97;
    ram_cell[     590] = 32'h0e72ae72;
    ram_cell[     591] = 32'h1c8cb27f;
    ram_cell[     592] = 32'hc8f03fba;
    ram_cell[     593] = 32'h64379927;
    ram_cell[     594] = 32'h0afd5a75;
    ram_cell[     595] = 32'h64b45aea;
    ram_cell[     596] = 32'h277e64fa;
    ram_cell[     597] = 32'h3d92f0cc;
    ram_cell[     598] = 32'h37ef9300;
    ram_cell[     599] = 32'h722b902b;
    ram_cell[     600] = 32'hf0c491d6;
    ram_cell[     601] = 32'h7f0fc0ae;
    ram_cell[     602] = 32'h42c18777;
    ram_cell[     603] = 32'hf22f9105;
    ram_cell[     604] = 32'h7d82fc0b;
    ram_cell[     605] = 32'h360aeaf6;
    ram_cell[     606] = 32'hf90af768;
    ram_cell[     607] = 32'ha00ae719;
    ram_cell[     608] = 32'hd880d792;
    ram_cell[     609] = 32'hb826751b;
    ram_cell[     610] = 32'he8d5fb98;
    ram_cell[     611] = 32'h35d97781;
    ram_cell[     612] = 32'he1558db0;
    ram_cell[     613] = 32'hb6c88dd1;
    ram_cell[     614] = 32'h3628eff4;
    ram_cell[     615] = 32'hac1e4e8e;
    ram_cell[     616] = 32'h77e50db4;
    ram_cell[     617] = 32'h14bd672f;
    ram_cell[     618] = 32'h7b5f8802;
    ram_cell[     619] = 32'heeec4472;
    ram_cell[     620] = 32'h8b6ae7cc;
    ram_cell[     621] = 32'hebbc7723;
    ram_cell[     622] = 32'hb104ba3a;
    ram_cell[     623] = 32'h0f562d23;
    ram_cell[     624] = 32'h8188d6a1;
    ram_cell[     625] = 32'h516240d8;
    ram_cell[     626] = 32'h53d502ed;
    ram_cell[     627] = 32'h003e9f34;
    ram_cell[     628] = 32'hb1ca5a45;
    ram_cell[     629] = 32'hda92d74d;
    ram_cell[     630] = 32'he8621ea5;
    ram_cell[     631] = 32'hcd0305c3;
    ram_cell[     632] = 32'hab88d345;
    ram_cell[     633] = 32'h068219be;
    ram_cell[     634] = 32'h78fb73d5;
    ram_cell[     635] = 32'haa3440f6;
    ram_cell[     636] = 32'hd8ef4401;
    ram_cell[     637] = 32'hde498b21;
    ram_cell[     638] = 32'h3058d12b;
    ram_cell[     639] = 32'h2457e052;
    ram_cell[     640] = 32'hd23bb014;
    ram_cell[     641] = 32'h64d7a3fe;
    ram_cell[     642] = 32'h2e76d331;
    ram_cell[     643] = 32'h2e580e02;
    ram_cell[     644] = 32'hffb3d641;
    ram_cell[     645] = 32'ha859bb81;
    ram_cell[     646] = 32'heac7b03e;
    ram_cell[     647] = 32'h83984f21;
    ram_cell[     648] = 32'h477489b0;
    ram_cell[     649] = 32'h680f93a0;
    ram_cell[     650] = 32'h7f77b488;
    ram_cell[     651] = 32'hcd3147b9;
    ram_cell[     652] = 32'haaae3578;
    ram_cell[     653] = 32'h1598d761;
    ram_cell[     654] = 32'h8cacc9f0;
    ram_cell[     655] = 32'h54a64374;
    ram_cell[     656] = 32'h973aed9a;
    ram_cell[     657] = 32'h14535fcf;
    ram_cell[     658] = 32'hfe3be79a;
    ram_cell[     659] = 32'h523ee6ec;
    ram_cell[     660] = 32'h6c0ed39b;
    ram_cell[     661] = 32'heb63601a;
    ram_cell[     662] = 32'hfede290b;
    ram_cell[     663] = 32'ha8bb70cc;
    ram_cell[     664] = 32'h2d6e3cb1;
    ram_cell[     665] = 32'hcd9d23f6;
    ram_cell[     666] = 32'hefcededa;
    ram_cell[     667] = 32'h9521c501;
    ram_cell[     668] = 32'h3638a7af;
    ram_cell[     669] = 32'hbe29c0a2;
    ram_cell[     670] = 32'h43341f73;
    ram_cell[     671] = 32'h1a3825e1;
    ram_cell[     672] = 32'h8b6230bf;
    ram_cell[     673] = 32'h9ebd2777;
    ram_cell[     674] = 32'hf2e4f67f;
    ram_cell[     675] = 32'h92c6210c;
    ram_cell[     676] = 32'h07ae6a12;
    ram_cell[     677] = 32'h19e22625;
    ram_cell[     678] = 32'hd3630831;
    ram_cell[     679] = 32'h418f6abb;
    ram_cell[     680] = 32'h73855714;
    ram_cell[     681] = 32'h3d40ba73;
    ram_cell[     682] = 32'h8c17f723;
    ram_cell[     683] = 32'h6a8eaaab;
    ram_cell[     684] = 32'h8771adb9;
    ram_cell[     685] = 32'hdaf6283f;
    ram_cell[     686] = 32'h4eded008;
    ram_cell[     687] = 32'hd0d26554;
    ram_cell[     688] = 32'h370055dd;
    ram_cell[     689] = 32'hba9431d7;
    ram_cell[     690] = 32'h15428e24;
    ram_cell[     691] = 32'h371246c6;
    ram_cell[     692] = 32'hc2d91316;
    ram_cell[     693] = 32'h6cb20d50;
    ram_cell[     694] = 32'h0618f349;
    ram_cell[     695] = 32'hdeac130a;
    ram_cell[     696] = 32'hf88fefcd;
    ram_cell[     697] = 32'h44c325b0;
    ram_cell[     698] = 32'hfae4f013;
    ram_cell[     699] = 32'h68fd1467;
    ram_cell[     700] = 32'h25046cd5;
    ram_cell[     701] = 32'h945847c9;
    ram_cell[     702] = 32'h2d50b1e6;
    ram_cell[     703] = 32'h33b7dd33;
    ram_cell[     704] = 32'hd896693e;
    ram_cell[     705] = 32'h5785f421;
    ram_cell[     706] = 32'hdbea1570;
    ram_cell[     707] = 32'h9eafb8cb;
    ram_cell[     708] = 32'he081e8d2;
    ram_cell[     709] = 32'h13b892f0;
    ram_cell[     710] = 32'hea52b3e8;
    ram_cell[     711] = 32'he5e1ed41;
    ram_cell[     712] = 32'h4bf89012;
    ram_cell[     713] = 32'h5bd0fc0f;
    ram_cell[     714] = 32'h0e4bdc21;
    ram_cell[     715] = 32'h080a0306;
    ram_cell[     716] = 32'hb087c51e;
    ram_cell[     717] = 32'h6a673d42;
    ram_cell[     718] = 32'h9d865c9d;
    ram_cell[     719] = 32'h5eff0d0b;
    ram_cell[     720] = 32'h05e018af;
    ram_cell[     721] = 32'h699f5583;
    ram_cell[     722] = 32'hd55b83f2;
    ram_cell[     723] = 32'h8fb2181d;
    ram_cell[     724] = 32'h7f900bf5;
    ram_cell[     725] = 32'h4fa2f869;
    ram_cell[     726] = 32'h89fa4e0f;
    ram_cell[     727] = 32'h3e58224b;
    ram_cell[     728] = 32'h3688aba0;
    ram_cell[     729] = 32'hd02a643a;
    ram_cell[     730] = 32'h4404f89f;
    ram_cell[     731] = 32'hc666177b;
    ram_cell[     732] = 32'ha668e141;
    ram_cell[     733] = 32'he58c846f;
    ram_cell[     734] = 32'hd1cfa2b2;
    ram_cell[     735] = 32'h3b4a4668;
    ram_cell[     736] = 32'h22860e2e;
    ram_cell[     737] = 32'h64e3a636;
    ram_cell[     738] = 32'h451e85ae;
    ram_cell[     739] = 32'h0f66d795;
    ram_cell[     740] = 32'hc6cf02bb;
    ram_cell[     741] = 32'h63ead421;
    ram_cell[     742] = 32'hb10e37fc;
    ram_cell[     743] = 32'had527114;
    ram_cell[     744] = 32'h0748624f;
    ram_cell[     745] = 32'h3a150d5f;
    ram_cell[     746] = 32'h8944c367;
    ram_cell[     747] = 32'h15c15a67;
    ram_cell[     748] = 32'h5fbb2d11;
    ram_cell[     749] = 32'h1b488cc6;
    ram_cell[     750] = 32'h920c166d;
    ram_cell[     751] = 32'h4208fa29;
    ram_cell[     752] = 32'h227f0ca3;
    ram_cell[     753] = 32'h66a1fd5c;
    ram_cell[     754] = 32'h3174ae7f;
    ram_cell[     755] = 32'haed67752;
    ram_cell[     756] = 32'hb51b2c76;
    ram_cell[     757] = 32'h4aecae31;
    ram_cell[     758] = 32'hbc1b98ee;
    ram_cell[     759] = 32'h562fc38e;
    ram_cell[     760] = 32'h968ea64c;
    ram_cell[     761] = 32'h39ce1808;
    ram_cell[     762] = 32'hfdc85e6c;
    ram_cell[     763] = 32'hdeceb6e9;
    ram_cell[     764] = 32'h22a86b7f;
    ram_cell[     765] = 32'h73186740;
    ram_cell[     766] = 32'h696bad77;
    ram_cell[     767] = 32'h27a01482;
end

endmodule
